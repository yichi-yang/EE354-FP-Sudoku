/*
File     : divider_top_with_single_step.v 
Author   : Gandhi Puvvada
Revision  : 1.2, 2.0, 3.0 (to suit Nexys 4)
Date : Feb 15, 2008, 10/14/08, 2/22/2010, 2/12/2012, 2/17/2020
*/

/*
 
 ******* Important difference to note *******
 In the divider_top.v for the divider simple, we had the Btn1 to serve as  
 the Start button and Btn0 to serve as the Ack button. Here, also we have 
 the same. This is different from the divider_with_debounce design. Here, we
 want to single-step the division while it is in compute state though we
 are running the core design at full 50MHz clock. We use Btn2 to single-step.
 ********************************************
 
*/
module sudoku_top        (   
        MemOE, MemWR, RamCS, QuadSpiFlashCS, // Disable the three memory chips

        ClkPort,                           // the 100 MHz incoming clock signal
        
        BtnL, BtnU, BtnD, BtnR,            // L = Prev, R = Next, U = Enter, D = Start
        BtnC,                              // the center button (this is our reset in most of our designs)
        Sw15, Sw3, Sw2, Sw1, Sw0,           // 5 switches
        Ld15, Ld6, Ld5, Ld4, Ld3, Ld2, Ld1, Ld0, // 8 LEDs
        An3, An2, An1, An0,                   // 4 anodes
        An7, An6, An5, An4,                // another 4 anodes (need turned off)
        Ca, Cb, Cc, Cd, Ce, Cf, Cg,        // 7 cathodes
        Dp                                 // Dot Point Cathode on SSDs
      );

     
                                
    /*  INPUTS */
    // Clock & Reset I/O
    input        ClkPort;    
    // Project Specific Inputs
    input        BtnL, BtnU, BtnD, BtnR, BtnC;    
    input        Sw15, Sw3, Sw2, Sw1, Sw0;
    
    
    /*  OUTPUTS */
    // Control signals on Memory chips     (to disable them)
    output      MemOE, MemWR, RamCS, QuadSpiFlashCS;
    // Project Specific Outputs
    // LEDs
    output      Ld0, Ld1, Ld2, Ld3, Ld4, Ld5, Ld6, Ld15;
    // SSD Outputs
    output      Cg, Cf, Ce, Cd, Cc, Cb, Ca, Dp;
    output      An0, An1, An2, An3;    
    output      An4, An5, An6, An7;

    
    /*  LOCAL SIGNALS */
    wire        Reset, ClkPort;
    wire        board_clk, sys_clk;
    wire [1:0]     ssdscan_clk;
    
    wire Prev, Next, Enter, Start, Clk;
    wire [3:0] InputValue;
    wire Init, Load, Forward, Check, Back, Disp, Fail;
    wire [3:0] Row, Col;
    wire [3:0] OutputValue, OutputAttempt;
    wire OutputFixed;


// to produce divided clock
    reg [26:0]    DIV_CLK;
// SSD (Seven Segment Display)
    reg [3:0]    SSD;
    wire [3:0]    SSD3, SSD2, SSD1, SSD0;
    reg [7:0]      SSD_CATHODES;
    
    
//------------    
// Disable the three memories so that they do not interfere with the rest of the design.
    assign {MemOE, MemWR, RamCS, QuadSpiFlashCS} = 4'b1111;
    
    
//------------
// CLOCK DIVISION

    // The clock division circuitary works like this:
    //
    // ClkPort ---> [BUFGP2] ---> board_clk
    // board_clk ---> [clock dividing counter] ---> DIV_CLK
    // DIV_CLK ---> [constant assignment] ---> sys_clk;
    
    BUFGP BUFGP1 (board_clk, ClkPort);     

// As the ClkPort signal travels throughout our design,
// it is necessary to provide global routing to this signal. 
// The BUFGPs buffer these input ports and connect them to the global 
// routing resources in the FPGA.

    // BUFGP BUFGP2 (Reset, BtnC); In the case of Spartan 3E (on Nexys-2 board), we were using BUFGP to provide global routing for the reset signal. But Spartan 6 (on Nexys-3) does not allow this.
    assign Reset = BtnC;
    
//------------
    // Our clock is too fast (100MHz) for SSD scanning
    // create a series of slower "divided" clocks
    // each successive bit is 1/2 frequency
  always @(posedge board_clk, posedge Reset)     
    begin                            
        if (Reset)
        DIV_CLK <= 0;
        else
        DIV_CLK <= DIV_CLK + 1'b1;
    end
//------------    
    // In this design, we run the core design at full 50MHz clock!
    assign    sys_clk = board_clk;
    // assign    sys_clk = DIV_CLK[25];


    //------------         

    assign InputValue = {Sw3, Sw2, Sw1, Sw0};
    
    // Unlike in the divider_simple, here we use one button BtnU to represent SCEN
    // Instantiate the debouncer    // module ee201_debouncer(CLK, RESET, PB, DPB, SCEN, MCEN, CCEN);
    // notice the "SCEN" is produced here and is sent into the divider core further below
ee201_debouncer #(.N_dc(25)) ee201_debouncer_1 
        (.CLK(sys_clk), .RESET(Reset), .PB(BtnU), .DPB( ), .SCEN( ), .MCEN(Enter), .CCEN( ));
ee201_debouncer #(.N_dc(25)) ee201_debouncer_2
        (.CLK(sys_clk), .RESET(Reset), .PB(BtnL), .DPB( ), .SCEN( ), .MCEN(Prev), .CCEN( ));
ee201_debouncer #(.N_dc(25)) ee201_debouncer_3
        (.CLK(sys_clk), .RESET(Reset), .PB(BtnR), .DPB( ), .SCEN( ), .MCEN(Next), .CCEN( ));
ee201_debouncer #(.N_dc(25)) ee201_debouncer_4
        (.CLK(sys_clk), .RESET(Reset), .PB(BtnD), .DPB( ), .SCEN(Start), .MCEN( ), .CCEN( ));
                            
                        
    // instantiate the core divider design. Note the .SCEN(SCEN)
SudokuSolver sudoku_1(.Prev(Prev), .Start(Start), .Next(Next), .Clk(sys_clk), .Reset(Reset),
                        .Enter(Enter), .OutputValue(OutputValue), .InputValue(InputValue),
                        .OutputAttempt(OutputAttempt), .Row(Row), .Col(Col), .Init(Init),
                        .Load(Load), .Forward(Forward), .Check(Check), .Back(Back),
                        .Disp(Disp), .Fail(Fail), .Single(Sw15), .OutputFixed(OutputFixed));

//------------
// OUTPUT: LEDS
    
    assign {Ld6, Ld5, Ld4, Ld3, Ld2, Ld1, Ld0} = {Init, Load, Forward, Check, Back, Disp, Fail};

    assign Ld15 = Sw15;

//------------
// SSD (Seven Segment Display)
    // reg [3:0]    SSD;
    // wire [3:0]    SSD3, SSD2, SSD1, SSD0;
    
    assign SSD3 = Row;
    assign SSD2 = Col;
    assign SSD1 = OutputValue;
    assign SSD0 = Check ? OutputAttempt : (Forward || Back || Disp) ? OutputFixed : InputValue;


    // need a scan clk for the seven segment display 
    
    // 100 MHz / 2^18 = 381.5 cycles/sec ==> frequency of DIV_CLK[17]
    // 100 MHz / 2^19 = 190.7 cycles/sec ==> frequency of DIV_CLK[18]
    // 100 MHz / 2^20 =  95.4 cycles/sec ==> frequency of DIV_CLK[19]
    
    // 381.5 cycles/sec (2.62 ms per digit) [which means all 4 digits are lit once every 10.5 ms (reciprocal of 95.4 cycles/sec)] works well.
    
    //                  --|  |--|  |--|  |--|  |--|  |--|  |--|  |--|  |   
    //                    |  |  |  |  |  |  |  |  |  |  |  |  |  |  |  | 
    //  DIV_CLK[17]       |__|  |__|  |__|  |__|  |__|  |__|  |__|  |__|
    //
    //               -----|     |-----|     |-----|     |-----|     |
    //                    |  0  |  1  |  0  |  1  |     |     |     |     
    //  DIV_CLK[18]       |_____|     |_____|     |_____|     |_____|
    //
    //         -----------|           |-----------|           |
    //                    |  0     0  |  1     1  |           |           
    //  DIV_CLK[19]       |___________|           |___________|
    //
    
    assign ssdscan_clk = DIV_CLK[19:18];

    assign An0    = !(~(ssdscan_clk[1]) && ~(ssdscan_clk[0]));  // when ssdscan_clk = 00
    assign An1    = !(~(ssdscan_clk[1]) &&  (ssdscan_clk[0]));  // when ssdscan_clk = 01
    assign An2    =  !((ssdscan_clk[1]) && ~(ssdscan_clk[0]));  // when ssdscan_clk = 10
    assign An3    =  !((ssdscan_clk[1]) &&  (ssdscan_clk[0]));  // when ssdscan_clk = 11
    assign {An7, An6, An5, An4} = 4'b1111;
    
    
    always @ (ssdscan_clk, SSD0, SSD1, SSD2, SSD3)
    begin : SSD_SCAN_OUT
        case (ssdscan_clk) 
                  2'b00: SSD = SSD0;
                  2'b01: SSD = SSD1;
                  2'b10: SSD = SSD2;
                  2'b11: SSD = SSD3;
        endcase 
    end

    // Following is Hex-to-SSD conversion
    always @ (SSD) 
    begin : HEX_TO_SSD
        case (SSD) // in this solution file the dot points are made to glow by making Dp = 0
            //                                                                abcdefg,Dp
            4'b0000: SSD_CATHODES = 8'b00000010; // 0
            4'b0001: SSD_CATHODES = 8'b10011110; // 1
            4'b0010: SSD_CATHODES = 8'b00100100; // 2
            4'b0011: SSD_CATHODES = 8'b00001100; // 3
            4'b0100: SSD_CATHODES = 8'b10011000; // 4
            4'b0101: SSD_CATHODES = 8'b01001000; // 5
            4'b0110: SSD_CATHODES = 8'b01000000; // 6
            4'b0111: SSD_CATHODES = 8'b00011110; // 7
            4'b1000: SSD_CATHODES = 8'b00000000; // 8
            4'b1001: SSD_CATHODES = 8'b00001000; // 9
            4'b1010: SSD_CATHODES = 8'b00010000; // A
            4'b1011: SSD_CATHODES = 8'b11000000; // B
            4'b1100: SSD_CATHODES = 8'b01100010; // C
            4'b1101: SSD_CATHODES = 8'b10000100; // D
            4'b1110: SSD_CATHODES = 8'b01100000; // E
            4'b1111: SSD_CATHODES = 8'b01110000; // F    
            default: SSD_CATHODES = 8'bXXXXXXXX; // default is not needed as we covered all cases
        endcase
    end    
    
    // reg [7:0]  SSD_CATHODES;
    assign {Ca, Cb, Cc, Cd, Ce, Cf, Cg, Dp} = {SSD_CATHODES[7:1], 1'b1};
    
endmodule
